//=====================================================================
// File   : sim_common.vh
// Brief  : Common simulation settings
//=====================================================================
`timescale 1ns/1ps

// System clock period for simulation (50 MHz -> 20 ns)
`define TCLK_NS 20